`timescale 1ns / 1ps
/////////////////////////////////////////////////////////
module lab5(
  input clk,
  input reset_n,
  input [3:0] usr_btn,
  output [3:0] usr_led,
  output LCD_RS,
  output LCD_RW,
  output LCD_E,
  output [3:0] LCD_D
);

// turn off all the LEDs
assign usr_led = 4'b0000;

wire btn_level, btn_pressed;
reg prev_btn_level;
reg [127:0] row_A = "Press BTN3 to   "; // Initialize the text of the first row. 
reg [127:0] row_B = "show a message.."; // Initialize the text of the second row.
//newly add
//reg [127:0] row_A;
//reg [127:0] row_B;
reg [15:0] fibo[0:24];
reg clockwise = 1;
integer i;
reg [7:0] index = 1;
reg [7:0] index_2 = 1;
reg [30:0] count = 0;

reg [7:0] line1[0:3];
reg [7:0] line2[0:3];

reg [7:0] num[0:1];
reg [7:0] ten[0:1];

initial begin
    fibo[0] = 16'h0000;
    fibo[1] = 16'h0001;
    for(i = 2;i < 25;i = i + 1)begin
        fibo[i] = fibo[i - 1] + fibo[i - 2];
    end
end

LCD_module lcd0(
  .clk(clk),
  .reset(~reset_n),
  .row_A(row_A),
  .row_B(row_B),
  .LCD_E(LCD_E),
  .LCD_RS(LCD_RS),
  .LCD_RW(LCD_RW),
  .LCD_D(LCD_D)
);
    
debounce btn_db0(
  .clk(clk),
  .btn_input(usr_btn[3]),
  .btn_output(btn_level)
);
    
always @(posedge clk) begin
  if (~reset_n)
    prev_btn_level <= 1;
  else
    prev_btn_level <= btn_level;
end

assign btn_pressed = (btn_level == 1 && prev_btn_level == 0);

always @(posedge clk)begin
    if(~reset_n)begin
        clockwise <= 1;
        index <= 1;
        index_2 <= 1;
    end
    else if(btn_pressed)begin
        clockwise <= ~clockwise;
    end
    
    count <= (count < 70000000)?count + 1:0;

        num[0] <= (index < 10)? index + 8'b00110000: (index % 10) + 8'b00110000;
        ten[0] <= (index < 10)? 8'b00110000: ((index < 20)?8'b00110001:8'b00110010);
        if(index < 25)begin
            num[1] <= ((index + 1) < 10)? (index + 1) + 8'b00110000: ((index + 1) % 10) + 8'b00110000;
            ten[1] <= (index + 1 < 10)? 8'b00110000: ((index + 1 < 20)?8'b00110001:8'b00110010);
        end
        else begin
            num[1] <= 8'b00110000;
            ten[1] <= 8'b00110000;
        end
        line1[0] <= (fibo[index - 1][15-:4] < 4'b1010)?{4'b0011,fibo[index - 1][15-:4] } : {4'b0100,(fibo[index - 1][15-:4] - 4'b1001) };
        line1[1] <= (fibo[index - 1][11-:4] < 4'b1010)?{4'b0011,fibo[index - 1][11-:4] } : {4'b0100,(fibo[index - 1][11-:4] - 4'b1001) };
        line1[2] <= (fibo[index - 1][7-:4] < 4'b1010)?{4'b0011,fibo[index - 1][7-:4] } : {4'b0100,(fibo[index - 1][7-:4] - 4'b1001) };
        line1[3] <= (fibo[index - 1][3:0] < 4'b1010)?{4'b0011,fibo[index - 1][3:0] } : {4'b0100,(fibo[index - 1][3:0] - 4'b1001) };
        //line1[0] <= (fibo[index_2 - 1][15-:4] < 4'b1010) ? {4'b0011,fibo[index_2 - 1][15-:4] } : {4'b0100,(fibo[index_2 - 1][15-:4] - 4'b1001) };
        //line1[1] <= (fibo[index_2 - 1][11-:4] < 4'b1010) ? {4'b0011,fibo[index_2 - 1][11-:4] } : {4'b0100,(fibo[index_2 - 1][11-:4] - 4'b1001) };
        //line1[2] <= (fibo[index_2 - 1][7-:4] < 4'b1010) ? {4'b0011,fibo[index_2 - 1][7-:4] } : {4'b0100,(fibo[index_2 - 1][7-:4] - 4'b1001) };
        //line1[3] <= (fibo[index_2 - 1][3:0] < 4'b1010) ? {4'b0011,fibo[index_2 - 1][3:0] } : {4'b0100,(fibo[index_2 - 1][3:0] - 4'b1001) };
        
        //line2[0] <= (fibo[ ((index < 8'b00011001)?index:0) ][15-:4] < 4'b1010)?{4'b0011,fibo[((index < 8'b00011001)?index:0)][15-:4] } : {4'b0100,(fibo[((index < 8'b00011001)?index:0)][15-:4] - 4'b1001) };
        //line2[1] <= (fibo[ ((index < 8'b00011001)?index:0) ][11-:4] < 4'b1010)?{4'b0011,fibo[((index < 8'b00011001)?index:0)][11-:4] } : {4'b0100,(fibo[((index < 8'b00011001)?index:0)][11-:4] - 4'b1001) };
        //line2[2] <= (fibo[ ((index < 8'b00011001)?index:0) ][7-:4] < 4'b1010)?{4'b0011,fibo[((index < 8'b00011001)?index:0)][7-:4] } : {4'b0100,(fibo[((index < 8'b00011001)?index:0)][7-:4] - 4'b1001) };
        //line2[3] <= (fibo[ ((index < 8'b00011001)?index:0) ][3:0] < 4'b1010)?{4'b0011,fibo[((index < 8'b00011001)?index:0)][3:0] } : {4'b0100,(fibo[((index < 8'b00011001)?index:0)][3:0] - 4'b1001) };
        //line2[0] <= (fibo[22][15-:4] < 4'b1010)?{4'b0011,fibo[22][15-:4] } : {4'b0100,(fibo[22][15-:4] - 4'b1001) };
        //line2[1] <= (fibo[22][11-:4] < 4'b1010)?{4'b0011,fibo[22][11-:4] } : {4'b0100,(fibo[22][11-:4] - 4'b1001) };
        //line2[2] <= (fibo[22][7-:4] < 4'b1010)?{4'b0011,fibo[22][7-:4] } : {4'b0100,(fibo[22][7-:4] - 4'b1001) };
        //line2[3] <= (fibo[22][3:0] < 4'b1010)?{4'b0011,fibo[22][3:0] } : {4'b0100,(fibo[22][3:0] - 4'b1001) };
        
        case(index)
            1 : begin
                line2[0] <= (fibo[1][15-:4] < 4'b1010)?{4'b0011,fibo[1][15-:4] } : {4'b0100,(fibo[1][15-:4] - 4'b1001) };
                line2[1] <= (fibo[1][11-:4] < 4'b1010)?{4'b0011,fibo[1][11-:4] } : {4'b0100,(fibo[1][11-:4] - 4'b1001) };
                line2[2] <= (fibo[1][7-:4] < 4'b1010)?{4'b0011,fibo[1][7-:4] } : {4'b0100,(fibo[1][7-:4] - 4'b1001) };
                line2[3] <= (fibo[1][3:0] < 4'b1010)?{4'b0011,fibo[1][3:0] } : {4'b0100,(fibo[1][3:0] - 4'b1001) };
            end
            2 : begin
                line2[0] <= (fibo[2][15-:4] < 4'b1010)?{4'b0011,fibo[2][15-:4] } : {4'b0100,(fibo[2][15-:4] - 4'b1001) };
                line2[1] <= (fibo[2][11-:4] < 4'b1010)?{4'b0011,fibo[2][11-:4] } : {4'b0100,(fibo[2][11-:4] - 4'b1001) };
                line2[2] <= (fibo[2][7-:4] < 4'b1010)?{4'b0011,fibo[2][7-:4] } : {4'b0100,(fibo[2][7-:4] - 4'b1001) };
                line2[3] <= (fibo[2][3:0] < 4'b1010)?{4'b0011,fibo[2][3:0] } : {4'b0100,(fibo[2][3:0] - 4'b1001) };
            end 
            3 : begin
                line2[0] <= (fibo[3][15-:4] < 4'b1010)?{4'b0011,fibo[3][15-:4] } : {4'b0100,(fibo[3][15-:4] - 4'b1001) };
                line2[1] <= (fibo[3][11-:4] < 4'b1010)?{4'b0011,fibo[3][11-:4] } : {4'b0100,(fibo[3][11-:4] - 4'b1001) };
                line2[2] <= (fibo[3][7-:4] < 4'b1010)?{4'b0011,fibo[3][7-:4] } : {4'b0100,(fibo[3][7-:4] - 4'b1001) };
                line2[3] <= (fibo[3][3:0] < 4'b1010)?{4'b0011,fibo[3][3:0] } : {4'b0100,(fibo[3][3:0] - 4'b1001) };
            end
            4 : begin
                line2[0] <= (fibo[4][15-:4] < 4'b1010)?{4'b0011,fibo[4][15-:4] } : {4'b0100,(fibo[4][15-:4] - 4'b1001) };
                line2[1] <= (fibo[4][11-:4] < 4'b1010)?{4'b0011,fibo[4][11-:4] } : {4'b0100,(fibo[4][11-:4] - 4'b1001) };
                line2[2] <= (fibo[4][7-:4] < 4'b1010)?{4'b0011,fibo[4][7-:4] } : {4'b0100,(fibo[4][7-:4] - 4'b1001) };
                line2[3] <= (fibo[4][3:0] < 4'b1010)?{4'b0011,fibo[4][3:0] } : {4'b0100,(fibo[4][3:0] - 4'b1001) };
            end
            5 : begin
                line2[0] <= (fibo[5][15-:4] < 4'b1010)?{4'b0011,fibo[5][15-:4] } : {4'b0100,(fibo[5][15-:4] - 4'b1001) };
                line2[1] <= (fibo[5][11-:4] < 4'b1010)?{4'b0011,fibo[5][11-:4] } : {4'b0100,(fibo[5][11-:4] - 4'b1001) };
                line2[2] <= (fibo[5][7-:4] < 4'b1010)?{4'b0011,fibo[5][7-:4] } : {4'b0100,(fibo[5][7-:4] - 4'b1001) };
                line2[3] <= (fibo[5][3:0] < 4'b1010)?{4'b0011,fibo[5][3:0] } : {4'b0100,(fibo[5][3:0] - 4'b1001) };
            end
            6 : begin
                line2[0] <= (fibo[6][15-:4] < 4'b1010)?{4'b0011,fibo[6][15-:4] } : {4'b0100,(fibo[6][15-:4] - 4'b1001) };
                line2[1] <= (fibo[6][11-:4] < 4'b1010)?{4'b0011,fibo[6][11-:4] } : {4'b0100,(fibo[6][11-:4] - 4'b1001) };
                line2[2] <= (fibo[6][7-:4] < 4'b1010)?{4'b0011,fibo[6][7-:4] } : {4'b0100,(fibo[6][7-:4] - 4'b1001) };
                line2[3] <= (fibo[6][3:0] < 4'b1010)?{4'b0011,fibo[6][3:0] } : {4'b0100,(fibo[6][3:0] - 4'b1001) };
            end
            7 : begin
                line2[0] <= (fibo[7][15-:4] < 4'b1010)?{4'b0011,fibo[7][15-:4] } : {4'b0100,(fibo[7][15-:4] - 4'b1001) };
                line2[1] <= (fibo[7][11-:4] < 4'b1010)?{4'b0011,fibo[7][11-:4] } : {4'b0100,(fibo[7][11-:4] - 4'b1001) };
                line2[2] <= (fibo[7][7-:4] < 4'b1010)?{4'b0011,fibo[7][7-:4] } : {4'b0100,(fibo[7][7-:4] - 4'b1001) };
                line2[3] <= (fibo[7][3:0] < 4'b1010)?{4'b0011,fibo[7][3:0] } : {4'b0100,(fibo[7][3:0] - 4'b1001) };
            end
            8 : begin
                line2[0] <= (fibo[8][15-:4] < 4'b1010)?{4'b0011,fibo[8][15-:4] } : {4'b0100,(fibo[8][15-:4] - 4'b1001) };
                line2[1] <= (fibo[8][11-:4] < 4'b1010)?{4'b0011,fibo[8][11-:4] } : {4'b0100,(fibo[8][11-:4] - 4'b1001) };
                line2[2] <= (fibo[8][7-:4] < 4'b1010)?{4'b0011,fibo[8][7-:4] } : {4'b0100,(fibo[8][7-:4] - 4'b1001) };
                line2[3] <= (fibo[8][3:0] < 4'b1010)?{4'b0011,fibo[8][3:0] } : {4'b0100,(fibo[8][3:0] - 4'b1001) };
            end
            9 : begin
                line2[0] <= (fibo[9][15-:4] < 4'b1010)?{4'b0011,fibo[9][15-:4] } : {4'b0100,(fibo[9][15-:4] - 4'b1001) };
                line2[1] <= (fibo[9][11-:4] < 4'b1010)?{4'b0011,fibo[9][11-:4] } : {4'b0100,(fibo[9][11-:4] - 4'b1001) };
                line2[2] <= (fibo[9][7-:4] < 4'b1010)?{4'b0011,fibo[9][7-:4] } : {4'b0100,(fibo[9][7-:4] - 4'b1001) };
                line2[3] <= (fibo[9][3:0] < 4'b1010)?{4'b0011,fibo[9][3:0] } : {4'b0100,(fibo[9][3:0] - 4'b1001) };
            end
            10 : begin
                line2[0] <= (fibo[10][15-:4] < 4'b1010)?{4'b0011,fibo[10][15-:4] } : {4'b0100,(fibo[10][15-:4] - 4'b1001) };
                line2[1] <= (fibo[10][11-:4] < 4'b1010)?{4'b0011,fibo[10][11-:4] } : {4'b0100,(fibo[10][11-:4] - 4'b1001) };
                line2[2] <= (fibo[10][7-:4] < 4'b1010)?{4'b0011,fibo[10][7-:4] } : {4'b0100,(fibo[10][7-:4] - 4'b1001) };
                line2[3] <= (fibo[10][3:0] < 4'b1010)?{4'b0011,fibo[10][3:0] } : {4'b0100,(fibo[10][3:0] - 4'b1001) };
            end
            11 : begin
                line2[0] <= (fibo[11][15-:4] < 4'b1010)?{4'b0011,fibo[11][15-:4] } : {4'b0100,(fibo[11][15-:4] - 4'b1001) };
                line2[1] <= (fibo[11][11-:4] < 4'b1010)?{4'b0011,fibo[11][11-:4] } : {4'b0100,(fibo[11][11-:4] - 4'b1001) };
                line2[2] <= (fibo[11][7-:4] < 4'b1010)?{4'b0011,fibo[11][7-:4] } : {4'b0100,(fibo[11][7-:4] - 4'b1001) };
                line2[3] <= (fibo[11][3:0] < 4'b1010)?{4'b0011,fibo[11][3:0] } : {4'b0100,(fibo[11][3:0] - 4'b1001) };
            end
            12 : begin
                line2[0] <= (fibo[12][15-:4] < 4'b1010)?{4'b0011,fibo[12][15-:4] } : {4'b0100,(fibo[12][15-:4] - 4'b1001) };
                line2[1] <= (fibo[12][11-:4] < 4'b1010)?{4'b0011,fibo[12][11-:4] } : {4'b0100,(fibo[12][11-:4] - 4'b1001) };
                line2[2] <= (fibo[12][7-:4] < 4'b1010)?{4'b0011,fibo[12][7-:4] } : {4'b0100,(fibo[12][7-:4] - 4'b1001) };
                line2[3] <= (fibo[12][3:0] < 4'b1010)?{4'b0011,fibo[12][3:0] } : {4'b0100,(fibo[12][3:0] - 4'b1001) };
            end
            13 : begin
                line2[0] <= (fibo[13][15-:4] < 4'b1010)?{4'b0011,fibo[13][15-:4] } : {4'b0100,(fibo[13][15-:4] - 4'b1001) };
                line2[1] <= (fibo[13][11-:4] < 4'b1010)?{4'b0011,fibo[13][11-:4] } : {4'b0100,(fibo[13][11-:4] - 4'b1001) };
                line2[2] <= (fibo[13][7-:4] < 4'b1010)?{4'b0011,fibo[13][7-:4] } : {4'b0100,(fibo[13][7-:4] - 4'b1001) };
                line2[3] <= (fibo[13][3:0] < 4'b1010)?{4'b0011,fibo[13][3:0] } : {4'b0100,(fibo[13][3:0] - 4'b1001) };
            end
            14 : begin
                line2[0] <= (fibo[14][15-:4] < 4'b1010)?{4'b0011,fibo[14][15-:4] } : {4'b0100,(fibo[14][15-:4] - 4'b1001) };
                line2[1] <= (fibo[14][11-:4] < 4'b1010)?{4'b0011,fibo[14][11-:4] } : {4'b0100,(fibo[14][11-:4] - 4'b1001) };
                line2[2] <= (fibo[14][7-:4] < 4'b1010)?{4'b0011,fibo[14][7-:4] } : {4'b0100,(fibo[14][7-:4] - 4'b1001) };
                line2[3] <= (fibo[14][3:0] < 4'b1010)?{4'b0011,fibo[14][3:0] } : {4'b0100,(fibo[14][3:0] - 4'b1001) };
            end
            15 : begin
                line2[0] <= (fibo[15][15-:4] < 4'b1010)?{4'b0011,fibo[15][15-:4] } : {4'b0100,(fibo[15][15-:4] - 4'b1001) };
                line2[1] <= (fibo[15][11-:4] < 4'b1010)?{4'b0011,fibo[15][11-:4] } : {4'b0100,(fibo[15][11-:4] - 4'b1001) };
                line2[2] <= (fibo[15][7-:4] < 4'b1010)?{4'b0011,fibo[15][7-:4] } : {4'b0100,(fibo[15][7-:4] - 4'b1001) };
                line2[3] <= (fibo[15][3:0] < 4'b1010)?{4'b0011,fibo[15][3:0] } : {4'b0100,(fibo[15][3:0] - 4'b1001) };
            end
            16 : begin
                line2[0] <= (fibo[16][15-:4] < 4'b1010)?{4'b0011,fibo[16][15-:4] } : {4'b0100,(fibo[16][15-:4] - 4'b1001) };
                line2[1] <= (fibo[16][11-:4] < 4'b1010)?{4'b0011,fibo[16][11-:4] } : {4'b0100,(fibo[16][11-:4] - 4'b1001) };
                line2[2] <= (fibo[16][7-:4] < 4'b1010)?{4'b0011,fibo[16][7-:4] } : {4'b0100,(fibo[16][7-:4] - 4'b1001) };
                line2[3] <= (fibo[16][3:0] < 4'b1010)?{4'b0011,fibo[16][3:0] } : {4'b0100,(fibo[16][3:0] - 4'b1001) };
            end
            17 : begin
                line2[0] <= (fibo[17][15-:4] < 4'b1010)?{4'b0011,fibo[17][15-:4] } : {4'b0100,(fibo[17][15-:4] - 4'b1001) };
                line2[1] <= (fibo[17][11-:4] < 4'b1010)?{4'b0011,fibo[17][11-:4] } : {4'b0100,(fibo[17][11-:4] - 4'b1001) };
                line2[2] <= (fibo[17][7-:4] < 4'b1010)?{4'b0011,fibo[17][7-:4] } : {4'b0100,(fibo[17][7-:4] - 4'b1001) };
                line2[3] <= (fibo[17][3:0] < 4'b1010)?{4'b0011,fibo[17][3:0] } : {4'b0100,(fibo[17][3:0] - 4'b1001) };
            end
            18 : begin
                line2[0] <= (fibo[18][15-:4] < 4'b1010)?{4'b0011,fibo[18][15-:4] } : {4'b0100,(fibo[18][15-:4] - 4'b1001) };
                line2[1] <= (fibo[18][11-:4] < 4'b1010)?{4'b0011,fibo[18][11-:4] } : {4'b0100,(fibo[18][11-:4] - 4'b1001) };
                line2[2] <= (fibo[18][7-:4] < 4'b1010)?{4'b0011,fibo[18][7-:4] } : {4'b0100,(fibo[18][7-:4] - 4'b1001) };
                line2[3] <= (fibo[18][3:0] < 4'b1010)?{4'b0011,fibo[18][3:0] } : {4'b0100,(fibo[18][3:0] - 4'b1001) };
            end
            19 : begin
                line2[0] <= (fibo[19][15-:4] < 4'b1010)?{4'b0011,fibo[19][15-:4] } : {4'b0100,(fibo[19][15-:4] - 4'b1001) };
                line2[1] <= (fibo[19][11-:4] < 4'b1010)?{4'b0011,fibo[19][11-:4] } : {4'b0100,(fibo[19][11-:4] - 4'b1001) };
                line2[2] <= (fibo[19][7-:4] < 4'b1010)?{4'b0011,fibo[19][7-:4] } : {4'b0100,(fibo[19][7-:4] - 4'b1001) };
                line2[3] <= (fibo[19][3:0] < 4'b1010)?{4'b0011,fibo[19][3:0] } : {4'b0100,(fibo[19][3:0] - 4'b1001) };
            end
            20 : begin
                line2[0] <= (fibo[20][15-:4] < 4'b1010)?{4'b0011,fibo[20][15-:4] } : {4'b0100,(fibo[20][15-:4] - 4'b1001) };
                line2[1] <= (fibo[20][11-:4] < 4'b1010)?{4'b0011,fibo[20][11-:4] } : {4'b0100,(fibo[20][11-:4] - 4'b1001) };
                line2[2] <= (fibo[20][7-:4] < 4'b1010)?{4'b0011,fibo[20][7-:4] } : {4'b0100,(fibo[20][7-:4] - 4'b1001) };
                line2[3] <= (fibo[20][3:0] < 4'b1010)?{4'b0011,fibo[20][3:0] } : {4'b0100,(fibo[20][3:0] - 4'b1001) };
            end
            21 : begin
                line2[0] <= (fibo[21][15-:4] < 4'b1010)?{4'b0011,fibo[21][15-:4] } : {4'b0100,(fibo[21][15-:4] - 4'b1001) };
                line2[1] <= (fibo[21][11-:4] < 4'b1010)?{4'b0011,fibo[21][11-:4] } : {4'b0100,(fibo[21][11-:4] - 4'b1001) };
                line2[2] <= (fibo[21][7-:4] < 4'b1010)?{4'b0011,fibo[21][7-:4] } : {4'b0100,(fibo[21][7-:4] - 4'b1001) };
                line2[3] <= (fibo[21][3:0] < 4'b1010)?{4'b0011,fibo[21][3:0] } : {4'b0100,(fibo[21][3:0] - 4'b1001) };
            end
            22 : begin
                line2[0] <= (fibo[22][15-:4] < 4'b1010)?{4'b0011,fibo[22][15-:4] } : {4'b0100,(fibo[22][15-:4] - 4'b1001) };
                line2[1] <= (fibo[22][11-:4] < 4'b1010)?{4'b0011,fibo[22][11-:4] } : {4'b0100,(fibo[22][11-:4] - 4'b1001) };
                line2[2] <= (fibo[22][7-:4] < 4'b1010)?{4'b0011,fibo[22][7-:4] } : {4'b0100,(fibo[22][7-:4] - 4'b1001) };
                line2[3] <= (fibo[22][3:0] < 4'b1010)?{4'b0011,fibo[22][3:0] } : {4'b0100,(fibo[22][3:0] - 4'b1001) };
            end
            23 : begin
                line2[0] <= (fibo[23][15-:4] < 4'b1010)?{4'b0011,fibo[23][15-:4] } : {4'b0100,(fibo[23][15-:4] - 4'b1001) };
                line2[1] <= (fibo[23][11-:4] < 4'b1010)?{4'b0011,fibo[23][11-:4] } : {4'b0100,(fibo[23][11-:4] - 4'b1001) };
                line2[2] <= (fibo[23][7-:4] < 4'b1010)?{4'b0011,fibo[23][7-:4] } : {4'b0100,(fibo[23][7-:4] - 4'b1001) };
                line2[3] <= (fibo[23][3:0] < 4'b1010)?{4'b0011,fibo[23][3:0] } : {4'b0100,(fibo[23][3:0] - 4'b1001) };
            end
            24 : begin
                line2[0] <= (fibo[24][15-:4] < 4'b1010)?{4'b0011,fibo[24][15-:4] } : {4'b0100,(fibo[24][15-:4] - 4'b1001) };
                line2[1] <= (fibo[24][11-:4] < 4'b1010)?{4'b0011,fibo[24][11-:4] } : {4'b0100,(fibo[24][11-:4] - 4'b1001) };
                line2[2] <= (fibo[24][7-:4] < 4'b1010)?{4'b0011,fibo[24][7-:4] } : {4'b0100,(fibo[24][7-:4] - 4'b1001) };
                line2[3] <= (fibo[24][3:0] < 4'b1010)?{4'b0011,fibo[24][3:0] } : {4'b0100,(fibo[24][3:0] - 4'b1001) };
            end
            25 : begin
                line2[0] <= (fibo[0][15-:4] < 4'b1010)?{4'b0011,fibo[0][15-:4] } : {4'b0100,(fibo[0][15-:4] - 4'b1001) };
                line2[1] <= (fibo[0][11-:4] < 4'b1010)?{4'b0011,fibo[0][11-:4] } : {4'b0100,(fibo[0][11-:4] - 4'b1001) };
                line2[2] <= (fibo[0][7-:4] < 4'b1010)?{4'b0011,fibo[0][7-:4] } : {4'b0100,(fibo[0][7-:4] - 4'b1001) };
                line2[3] <= (fibo[0][3:0] < 4'b1010)?{4'b0011,fibo[0][3:0] } : {4'b0100,(fibo[0][3:0] - 4'b1001) };
            end
            default : begin
                line2[0] <= (fibo[0][15-:4] < 4'b1010)?{4'b0011,fibo[0][15-:4] } : {4'b0100,(fibo[0][15-:4] - 4'b1001) };
                line2[1] <= (fibo[0][11-:4] < 4'b1010)?{4'b0011,fibo[0][11-:4] } : {4'b0100,(fibo[0][11-:4] - 4'b1001) };
                line2[2] <= (fibo[0][7-:4] < 4'b1010)?{4'b0011,fibo[0][7-:4] } : {4'b0100,(fibo[0][7-:4] - 4'b1001) };
                line2[3] <= (fibo[0][3:0] < 4'b1010)?{4'b0011,fibo[0][3:0] } : {4'b0100,(fibo[0][3:0] - 4'b1001) };
            end
            
        endcase

   
    if(count == 69999999)begin
        row_A <= {"Fibo #",ten[0],num[0]," is ",line1[0],line1[1],line1[2],line1[3]};
        row_B <= {"Fibo #",ten[1],num[1]," is ",line2[0],line2[1],line2[2],line2[3]};
        if(clockwise == 1)begin
            index <= (index < 25)?index + 1:1;
            index_2 <= (index_2 < 25)?index_2 + 1:1;
        end
        else if(clockwise == 0)begin
            index <= (index > 1)?index - 1:25;
            index_2 <= (index_2 > 1)?index_2 - 1:25;
        end
    end
end

endmodule

module debounce(
    input clk,
    input btn_input,
    output btn_output
    );
    assign btn_output = btn_input;
endmodule
